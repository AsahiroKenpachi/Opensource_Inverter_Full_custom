magic
tech sky130A
timestamp 1707906826
<< nwell >>
rect -150 -100 150 305
<< nmos >>
rect -10 -270 5 -170
<< pmos >>
rect -10 -50 5 150
<< ndiff >>
rect -50 -180 -10 -170
rect -50 -260 -45 -180
rect -25 -260 -10 -180
rect -50 -270 -10 -260
rect 5 -180 50 -170
rect 5 -260 20 -180
rect 40 -260 50 -180
rect 5 -270 50 -260
<< pdiff >>
rect -55 140 -10 150
rect -55 -40 -45 140
rect -25 -40 -10 140
rect -55 -50 -10 -40
rect 5 140 50 150
rect 5 -40 20 140
rect 40 -40 50 140
rect 5 -50 50 -40
<< ndiffc >>
rect -45 -260 -25 -180
rect 20 -260 40 -180
<< pdiffc >>
rect -45 -40 -25 140
rect 20 -40 40 140
<< psubdiff >>
rect -50 -340 50 -330
rect -50 -360 -30 -340
rect 30 -360 50 -340
rect -50 -370 50 -360
<< nsubdiff >>
rect -60 275 50 285
rect -60 255 -30 275
rect 30 255 50 275
rect -60 245 50 255
<< psubdiffcont >>
rect -30 -360 30 -340
<< nsubdiffcont >>
rect -30 255 30 275
<< poly >>
rect -10 150 5 200
rect -10 -105 5 -50
rect -75 -115 5 -105
rect -75 -140 -70 -115
rect -40 -140 5 -115
rect -75 -150 5 -140
rect 65 -115 115 -105
rect 65 -140 75 -115
rect 105 -140 115 -115
rect 65 -150 115 -140
rect -10 -170 5 -150
rect -10 -310 5 -270
<< polycont >>
rect -70 -140 -40 -115
rect 75 -140 105 -115
<< locali >>
rect -60 275 50 285
rect -60 255 -30 275
rect 30 255 50 275
rect -60 245 50 255
rect -55 150 -25 245
rect -55 140 -15 150
rect -55 -40 -45 140
rect -25 -40 -15 140
rect -55 -50 -15 -40
rect 10 140 50 150
rect 10 -40 20 140
rect 40 -40 50 140
rect 10 -50 50 -40
rect 15 -105 45 -50
rect -75 -115 -25 -105
rect -75 -140 -70 -115
rect -40 -140 -25 -115
rect -75 -150 -25 -140
rect 15 -115 115 -105
rect 15 -140 75 -115
rect 105 -140 115 -115
rect 15 -150 115 -140
rect 15 -170 45 -150
rect -50 -180 -15 -170
rect -50 -260 -45 -180
rect -25 -260 -15 -180
rect -50 -270 -15 -260
rect 10 -180 50 -170
rect 10 -260 20 -180
rect 40 -260 50 -180
rect 10 -270 50 -260
rect -45 -330 -20 -270
rect -50 -340 50 -330
rect -50 -360 -30 -340
rect 30 -360 50 -340
rect -50 -370 50 -360
<< viali >>
rect -25 255 20 275
rect -70 -140 -40 -115
rect 75 -140 105 -115
rect -15 -360 10 -340
<< metal1 >>
rect -185 275 215 285
rect -185 255 -25 275
rect 20 255 215 275
rect -185 245 215 255
rect -185 -115 -25 -105
rect -185 -140 -70 -115
rect -40 -140 -25 -115
rect -185 -150 -25 -140
rect 15 -115 265 -105
rect 15 -140 75 -115
rect 105 -140 265 -115
rect 15 -150 265 -140
rect -200 -340 195 -330
rect -200 -360 -15 -340
rect 10 -360 195 -340
rect -200 -375 195 -360
<< labels >>
rlabel metal1 263 -123 263 -123 7 vout
port 2 w
rlabel metal1 -181 -124 -181 -124 1 vin
port 3 n
rlabel metal1 194 -353 194 -353 1 gnd
port 4 n
rlabel metal1 206 271 206 271 1 v1
port 1 n
<< end >>
